//==================================================================================================
//  Note:          Use only for teaching materials of IC Design Lab, NTHU.
//  Copyright: (c) 2025 Vision Circuits and Systems Lab, NTHU, Taiwan. ALL Rights Reserved.
//==================================================================================================

module enigma(clk, srst_n, load, encrypt, crypt_mode, table_idx, code_in, code_out, code_valid);
input clk;         // clock 
input srst_n;      // synchronous reset (active low)
input load;        // load control signal (level sensitive). 0/1: inactive/active
input encrypt;     // encrypt control signal (level sensitive). 0/1: inactive/active
input crypt_mode;  // 0: encrypt; 1:decrypt;
input [2-1:0] table_idx; // table_idx indicates which rotor to be loaded 
						             // 2'b00: rotorA
						             // 2'b01: plugboard
						             // 2'b10: rotorB
input [6-1:0] code_in;	// When load is active, then code_in is input of rotors. 
						// When encrypy is active, then code_in is input of code words.
output reg [6-1:0] code_out;   // encrypted code word
output reg code_valid;         // 0: non-valid code_out; 1: valid code_out 

// ======== Declarations ======== //

wire XOR_whitening_en;
wire [5:0] XOR_whitening_in;
wire [5:0] XOR_whitening_out;
wire XOR_whitening_out_valid;

wire [5:0] rotorA_ls_count, rotorA_for_dout;
wire rotorA_for_out_valid;
wire rotorA_we;

wire [5:0] for_bit_sw_out, inv_bit_sw_out;

wire [5:0] rotorA_inv_dout;
wire rotorA_inv_out_valid;

reg load_ff, encrypt_ff, crypt_mode_ff;
reg [1:0] table_idx_ff;
reg [5:0] code_in_ff;

wire [5:0] rotorB_for_din, rotorB_for_dout;
wire [5:0] rotorB_inv_din, rotorB_inv_dout;
wire rotorB_for_in_valid, rotorB_inv_in_valid;
wire rotorB_for_out_valid, rotorB_inv_out_valid;

wire bit_sw_inv_out_valid, bit_sw_inv_in_valid;

// ======== Input ff ========== //


always @ (posedge clk) begin
  {load_ff, encrypt_ff, crypt_mode_ff, table_idx_ff, code_in_ff} <= {load, encrypt, crypt_mode, table_idx, code_in};
end


// ============ Plugboard ============= //

wire [5:0] plugboard_for_din, plugboard_inv_din; 
wire [5:0] plugboard_for_dout, plugboard_inv_dout;
wire plugboard_for_out_valid, plugboard_inv_out_valid;

assign plugboard_for_din = code_in_ff;
assign plugboard_inv_din = rotorA_inv_dout;

plugboard U_plugboard(
	.clk(clk),
	.srst_n(srst_n),
	.plugboard_for_din(plugboard_for_din), // = code_in_ff
	.plugboard_inv_din(plugboard_inv_din), // from rotorA
	.plugboard_for_dout(plugboard_for_dout),
	.plugboard_inv_dout(plugboard_inv_dout),
	.table_idx_ff(table_idx_ff),
	.load_ff(load_ff),
	.encrypt_ff(encrypt_ff),
	.plugboard_inv_in_valid(rotorA_inv_out_valid),
	.plugboard_for_out_valid(plugboard_for_out_valid),
	.plugboard_inv_out_valid(plugboard_inv_out_valid)
);



// ======== Rotor A (forward)========== //

rotorA_forward U_rotorA_forward(
  .clk(clk),
  .srst_n(srst_n),
  .rotorA_for_din(plugboard_for_dout), // write input (=code_in_ff in part123)
  .code_in_ff(code_in_ff),
  .table_idx_ff(table_idx_ff),
  .crypt_mode_ff(crypt_mode_ff),
  .encrypt_ff(plugboard_for_out_valid),
  .load_ff(load_ff),
  .inverse_path_LSB(inv_bit_sw_out[1:0]), // the least significant 2-bit of the input of the inverse pass
  .rotorA_for_dout(rotorA_for_dout), // read output
  .rotorA_ls_count(rotorA_ls_count), // the left shift count
  .rotorA_for_out_valid(rotorA_for_out_valid),
  .rotorA_we(rotorA_we)
);

// ========= Bit switching ========= //
//reg [5:0] rotorB_for_din_ff, rotorB_inv_dout_ff;

wire [5:0] inv_text_in;
assign inv_text_in = rotorB_inv_dout;
assign bit_sw_inv_in_valid = rotorB_inv_out_valid;

bit_sw U_bit_sw(
	.clk(clk),
  .srst_n(srst_n),
	.for_text_in(rotorA_for_dout),
	.inv_text_in(inv_text_in),
	.crypt_mode_ff(crypt_mode_ff),
	.sw_enable(rotorA_for_out_valid),
	.for_text_out(for_bit_sw_out),
	.inv_text_out(inv_bit_sw_out),
  .bit_sw_inv_in_valid(bit_sw_inv_in_valid),
  .bit_sw_inv_out_valid(bit_sw_inv_out_valid)
);

// ============ rotorB ============= //


/*
always @ (posedge clk) begin
  rotorB_for_din_ff <= rotorB_for_din;
  rotorB_inv_dout_ff <= rotorB_inv_dout;
end
*/

assign rotorB_for_din = for_bit_sw_out;
assign rotorB_inv_din = XOR_whitening_out;
assign rotorB_for_in_valid = rotorA_for_out_valid; // rotorA, bit sw, rotorB in same cycle
assign rotorB_inv_in_valid = XOR_whitening_out_valid;

rotorB U_rotorB(
	.clk(clk),
	.rotorB_for_din(rotorB_for_din), 
	.rotorB_inv_din(rotorB_inv_din),
	.rotorB_for_dout(rotorB_for_dout),
	.rotorB_inv_dout(rotorB_inv_dout),

	// control signals
	.rotorB_for_in_valid(rotorB_for_in_valid),
	.rotorB_inv_in_valid(rotorB_inv_in_valid),
	.code_in_ff(code_in_ff),
	.table_idx_ff(table_idx_ff),
	.crypt_mode_ff(crypt_mode_ff),
	.load_ff(load_ff),

	// output control signals
	.rotorB_for_out_valid(rotorB_for_out_valid),
	.rotorB_inv_out_valid(rotorB_inv_out_valid)
);

// ========= XOR Whitening ========= //

assign XOR_whitening_en = rotorB_for_out_valid;
assign XOR_whitening_in = rotorB_for_dout;

XOR_whitening U_XOR_whitening(
	.clk(clk),
	.srst_n(srst_n),
	.XOR_whitening_en(XOR_whitening_en),
	.XOR_whitening_in(XOR_whitening_in),
	.XOR_whitening_out(XOR_whitening_out),
	.XOR_whitening_out_valid(XOR_whitening_out_valid)
);

// ======== Rotor A (inverse)========== //
rotorA_inverse U_rotorA_inverse(
	.clk(clk),
	.srst_n(srst_n),
	.rotorA_inv_din(inv_bit_sw_out), // write input (=code_in_ff in part123)
	.rotorA_ls_count(rotorA_ls_count), // the left shift count
	.code_in_ff(code_in_ff),
	.rotorA_we(rotorA_we), // rotorA must share same we
	.rotorA_inv_dout(rotorA_inv_dout), // read output
	.rotorA_inv_in_valid(bit_sw_inv_out_valid),
	.rotorA_inv_out_valid(rotorA_inv_out_valid)
);

// ============ Final result =============== //

always @ (posedge clk) begin
  code_out    <= plugboard_inv_dout;
  code_valid  <= plugboard_inv_out_valid;
end

endmodule

//==============================================================//
//======================= Modules ==============================//
//==============================================================//

module sram64x6 (
  input        clk,
  input        we,    // write enable (1:write, 0:read)
  input  [5:0] addr, 
  input  [5:0] din,
  output [5:0] dout
);
  reg [5:0] mem [0:63];
  //reg [5:0] addr_r;

  always @(posedge clk) begin
    if (we) mem[addr] <= din;
    //addr_r <= addr;
  end
  assign dout = mem[addr];

endmodule

module sram64x6_rotorA_for (
  input        clk,
  input        load,    // load enable
  input  [5:0] addr, 
  input  [5:0] din,
  output [5:0] dout
);
  reg [5:0] mem [0:63];
  //reg [5:0] addr_r;
  integer i;

  always @(posedge clk) begin
    if (load) begin
		mem[63] <= din;
		for (i=0; i<63; i=i+1)
			mem[i] <= mem[i+1];
	end
  end
  assign dout = mem[addr];

endmodule


module XOR_whitening(
	input clk,
	input srst_n,
  input XOR_whitening_en,
  input [5:0] XOR_whitening_in,
	output [5:0] XOR_whitening_out,
  output XOR_whitening_out_valid
);

reg [5:0] state, state_next;

always @* begin
  if (XOR_whitening_en) state_next = {state[4:0], state[4]^state[5]};
  else state_next = state;
end

always @ (posedge clk) begin
  if (~srst_n) state <= 6'b000001;
  else state <= state_next;
end

/*
always @ (posedge clk) begin
  XOR_whitening_out <= XOR_whitening_in ^ state;
  XOR_whitening_out_valid <= XOR_whitening_en;
end
*/

assign  XOR_whitening_out = XOR_whitening_in ^ state;
assign  XOR_whitening_out_valid = XOR_whitening_en;

endmodule




module rotorA_forward (
  input clk,
  input srst_n,
  input [5:0] rotorA_for_din, // read request (=code_in_ff in part123)
  input [5:0] code_in_ff,
  input [1:0] table_idx_ff,
  input crypt_mode_ff,
  input encrypt_ff,
  input load_ff,
  input [1:0] inverse_path_LSB, // the least significant 2-bit of the input of the inverse pass
  output [5:0] rotorA_for_dout, // read output
  output reg [5:0] rotorA_ls_count, // the left shift count
  output reg rotorA_for_out_valid,
  output reg rotorA_we // rotorA must share same we
);



reg [5:0] rotorA_ls_count_next; // the left shift count
reg [5:0] rotorA_addr_for;
reg [5:0] rotorA_addr_for_next;
reg  rotorA_we_next;


// module connection
sram64x6_rotorA_for U_rotorA_forward_buffer(
  .clk(clk),
  .load(rotorA_we_next),
  .addr(rotorA_addr_for), 
  .din(code_in_ff),
  .dout(rotorA_for_dout)
);

// write enable
always @*
 rotorA_we_next = (table_idx_ff == 2'b00 && load_ff == 1'b1);


// we have to know which cycles have a valid rotor output
always @ (posedge clk) begin
  rotorA_for_out_valid <= encrypt_ff;
end


// rotor A left shift count
always @ * begin
	if (rotorA_we_next) rotorA_ls_count_next = rotorA_ls_count + 1;
	else if (rotorA_for_out_valid) rotorA_ls_count_next = (crypt_mode_ff) ? rotorA_ls_count + inverse_path_LSB : rotorA_ls_count + rotorA_for_dout[1:0]; // 0: encrypt; 1:decrypt;
  else rotorA_ls_count_next = rotorA_ls_count;
end



// address
always @ * begin
  if (encrypt_ff) begin // when encrypting
    rotorA_addr_for_next = rotorA_for_din + rotorA_ls_count_next;
  end
  else begin   // when loading rotorA (or maybe other parts)
    rotorA_addr_for_next = rotorA_ls_count;
  end
end

// ======================

// rotorA table's data FF
always @ (posedge clk) begin
  rotorA_we <= rotorA_we_next;
end

// table's address & ls_count FF
always @ (posedge clk) begin
	if (~srst_n) begin
		rotorA_ls_count <= 6'd0;
		rotorA_addr_for	<= 6'd0;
	end
	else begin
		rotorA_ls_count <= rotorA_ls_count_next;
		rotorA_addr_for	<= rotorA_addr_for_next;
	end
end


endmodule


module rotorA_inverse (
  input clk,
  input srst_n,
  input [5:0] rotorA_inv_din, 
  input  [5:0] rotorA_ls_count, // the left shift count
  input rotorA_we, // rotorA must share same we
  input [5:0] code_in_ff,
  output [5:0] rotorA_inv_dout, // read output

  input rotorA_inv_in_valid,
  output reg rotorA_inv_out_valid
);

reg [5:0]  rotorA_addr_inv, rotorA_din_inv;
reg [5:0] rotorA_addr_inv_next, rotorA_din_inv_next;
wire [5:0] rotorA_inv_sram_dout;

// module connection
sram64x6 U_rotorA_inverse_buffer(
  .clk(clk),
  .we(rotorA_we),
  .addr(rotorA_addr_inv), 
  .din(rotorA_din_inv),
  .dout(rotorA_inv_sram_dout)
);

// rotorA din
always @ * begin
    rotorA_din_inv_next = rotorA_ls_count;
end

// address
always @ * begin
  if (rotorA_inv_in_valid) rotorA_addr_inv_next = rotorA_inv_din;
  else rotorA_addr_inv_next = code_in_ff;
end

// current left shift count need to be add to result
reg [5:0] ls_count_buffer, ls_count_buffer_next;
wire [5:0] rotorA_inv_sram_dout_fixed;

always @ (posedge clk) begin
  ls_count_buffer <= rotorA_ls_count;
  rotorA_inv_out_valid <= rotorA_inv_in_valid;
end

assign rotorA_inv_dout = rotorA_inv_sram_dout - ls_count_buffer;


// rotorA table's data FF
always @ (posedge clk) begin
	rotorA_din_inv 	<= rotorA_din_inv_next;
end

// table's address & ls_count FF
always @ (posedge clk) begin
	if (~srst_n) begin
		rotorA_addr_inv	<= 6'd0;
	end
	else begin
		rotorA_addr_inv	<= rotorA_addr_inv_next;
	end
end

endmodule

module bit_sw(
	input clk,
	input srst_n,
	input [5:0] for_text_in,
	input [5:0] inv_text_in,
	input crypt_mode_ff,
	input sw_enable,
	output reg [5:0] for_text_out,
	output reg [5:0] inv_text_out,
  input bit_sw_inv_in_valid, 
  output bit_sw_inv_out_valid
);

reg [1:0] mode, mode_next;

assign bit_sw_inv_out_valid = bit_sw_inv_in_valid;

always @ * begin
	if (sw_enable) mode_next = (crypt_mode_ff) ? inv_text_in[1:0] : for_text_out[1:0];// 0: encrypt; 1:decrypt;
	else mode_next = mode;
end

always @* begin
	case(mode)
		2'b00: for_text_out = ~for_text_in;
		2'b01: for_text_out = {for_text_in[0], for_text_in[1], for_text_in[2], for_text_in[3], for_text_in[4], for_text_in[5]};
		2'b10: for_text_out = {for_text_in[4], for_text_in[5], for_text_in[2], for_text_in[3], for_text_in[0], for_text_in[1]};
		2'b11: for_text_out = {for_text_in[2], for_text_in[1], for_text_in[0], for_text_in[5], for_text_in[4], for_text_in[3]};
	endcase
end

always @* begin
	case(mode)
		2'b00: inv_text_out = ~inv_text_in;
		2'b01: inv_text_out = {inv_text_in[0], inv_text_in[1], inv_text_in[2], inv_text_in[3], inv_text_in[4], inv_text_in[5]};
		2'b10: inv_text_out = {inv_text_in[4], inv_text_in[5], inv_text_in[2], inv_text_in[3], inv_text_in[0], inv_text_in[1]};
		2'b11: inv_text_out = {inv_text_in[2], inv_text_in[1], inv_text_in[0], inv_text_in[5], inv_text_in[4], inv_text_in[3]};
	endcase
end

always @ (posedge clk) begin
	if (~srst_n) mode <= 0;
	else mode <= mode_next;
end

endmodule




module plugboard (
	input clk,
	input srst_n,
	input [5:0] plugboard_for_din, // = code_in_ff
	input [5:0] plugboard_inv_din, // from rotorA
	output [5:0] plugboard_for_dout,
	output [5:0] plugboard_inv_dout,

	input [1:0] table_idx_ff,
	input load_ff,
	input encrypt_ff,

	input plugboard_inv_in_valid,
	output reg plugboard_for_out_valid,
	output reg plugboard_inv_out_valid
);
// 2 cycles delay
// plugboard_for_din GET THE CORRESPONDING OUTPUT RESPONSE plugboard_for_dout AFTER 2 CYCLES

// 2 cycles read delay for inv too, TODO (may be reduce to 1 delay for better performance ?)

// ======== Declaration ========= //
reg state, state_next;
reg plugboard_we_next, plugboard_we, plugboard_we_ff;
//reg [5:0] plugboard_for_addr, plugboard_for_addr_next;
wire [5:0] plugboard_for_addr;
reg [5:0]  plugboard_inv_addr, plugboard_inv_addr_next;
//reg [5:0] plugboard_sram_din, plugboard_sram_din_next;
wire [5:0] plugboard_sram_din;
reg [17:0] temp;
reg plugboard_for_out_valid_beforeff;
reg plugboard_inv_out_valid_beforeff;

// module connection
sram2r1w_64x6 U_plugboard(
  .clk(clk),
  .srst_n(srst_n),
  .we(plugboard_we_ff),
  .addr_for(plugboard_for_addr), 
  .addr_inv(plugboard_inv_addr),
  .din(plugboard_sram_din),
  .dout_for(plugboard_for_dout),
  .dout_inv(plugboard_inv_dout)
);

// ============================== //

localparam CYCLE1 = 1'b0;
localparam CYCLE2 = 1'b1;

// write enable
always @*
	plugboard_we_next = (table_idx_ff == 2'b01 && load_ff == 1'b1);

// state control
always @* begin
	if (plugboard_we_ff) state_next = ~state;
	else state_next = CYCLE2; // addr = temp[5:0] (delay only 1 cycle)
end

// temp buffer (keep left shifting)
always @ (posedge clk) begin
	temp <= {temp[11:0], plugboard_for_din};
end

// cycle 1 : temp[17:0] <= {6'd?, 6'd?, in_cycle1[5:0]};
// cycle 2 : temp[17:0] <= {6'd?, in_cycle1[5:0], in_cycle2[5:0]};
// cycle 3 : temp[17:0] <= {in_cycle1[5:0], in_cycle2[5:0], in_cycle3[5:0]};
// cycle 4 : temp[17:0] <= {in_cycle2[5:0], in_cycle3[5:0], in_cycle4[5:0]};
	// addr = in_cycle1, data = in_cycle2;
	// addr = in_cycle2, data = in_cycle1;
	// CYCLE1 : addr = temp[17:12], data = temp[11:6];
	// CYCLE2 : addr = temp[5:0], data = temp[11:6];
	// first write start in cycle2
	// to minimize the delay, encrypt/decrypt in CYCLE2

// sram_din & addr_for control
assign plugboard_sram_din = temp[11:6];
assign plugboard_for_addr = state == CYCLE1 ? temp[17:12] : temp[5:0];

// addr_inv control
always @ * begin
	plugboard_inv_addr_next = plugboard_inv_din;
end



always @ (posedge clk) begin
	plugboard_we		<= plugboard_we_next;
	plugboard_we_ff		<= plugboard_we;
	state				<= state_next;
	//plugboard_sram_din 	<= plugboard_sram_din_next;
	plugboard_inv_addr					<= plugboard_inv_addr_next;
	//plugboard_inv_out_valid_beforeff	<= plugboard_inv_in_valid;
	//plugboard_inv_out_valid 			<= plugboard_inv_out_valid_beforeff;
	plugboard_inv_out_valid 			<= plugboard_inv_in_valid;
	plugboard_for_out_valid_beforeff 	<= encrypt_ff;
	plugboard_for_out_valid 			<= plugboard_for_out_valid_beforeff;
end

endmodule


module sram2r1w_64x6 (
  input        clk,
  input 	   srst_n,
  input        we,    			// write enable (1:write, 0:read)
  input  [5:0] addr_for, 		// forward address
  input  [5:0] addr_inv, 		// inverse address
  input  [5:0] din,				// input write data
  output reg [5:0] dout_for, 	// forward dout
  output [5:0] dout_inv 	// inverse dout
);
  reg [5:0] mem [0:63];
  integer i;

  always @(posedge clk) begin
	dout_for	<= mem[addr_for];
  end

  always @ (posedge clk) begin
	if (~srst_n) begin
		for(i=0; i<64; i=i+1) mem[i] <= i;
	end
	else if (we) mem[addr_for] <= din;
  end

  assign dout_inv = mem[addr_inv];

endmodule

module rotorB (
	input clk,
	input [5:0] rotorB_for_din, // read request (=code_in_ff in part123)
	input [5:0] rotorB_inv_din,
	output [5:0] rotorB_for_dout,
	output [5:0] rotorB_inv_dout,

	// control signals
	input rotorB_for_in_valid,
	input rotorB_inv_in_valid,
	input [5:0] code_in_ff,
	input [1:0] table_idx_ff,
	input crypt_mode_ff,
	input load_ff,

	// output control signals
	output rotorB_for_out_valid,
	output rotorB_inv_out_valid
);

wire load_sram; // load the 64 data
wire [1:0] rot_mode; // the stage1 rotor mode

// TODO simplfied : table_idx_ff[1] == 1;
assign load_sram = (table_idx_ff == 2'b10) && load_ff;
assign rot_mode = (crypt_mode_ff) ? rotorB_inv_din[1:0] : rotorB_for_dout[1:0] ;

sram64x6_rotorB U_sram64x6_rotorB(
  .clk(clk),
  .load(load_sram),    // load enable

  .rotorB_sram_din(code_in_ff),
  .rotorB_for_addr(rotorB_for_din), // input address
  .rotorB_inv_din(rotorB_inv_din), // input data

  .rotorB_for_dout(rotorB_for_dout),	//output data
  .rotorB_inv_dout(rotorB_inv_dout), // output address

  .rot_mode(rot_mode),
  .rotorB_in_valid(rotorB_for_in_valid)
);

assign rotorB_for_out_valid = rotorB_for_in_valid;
assign rotorB_inv_out_valid = rotorB_inv_in_valid;



endmodule


module sram64x6_rotorB (
  input        clk,
  input        load,    // load enable

  input  [5:0] rotorB_sram_din,
  input  [5:0] rotorB_for_addr, // input address
  input  [5:0] rotorB_inv_din, // input data

  output [5:0] rotorB_for_dout,	//output data
  output reg [5:0] rotorB_inv_dout, // output address

  input [1:0] rot_mode,
  input rotorB_in_valid
);

reg [5:0] mem [0:63];
//reg [5:0] addr_r;
integer i;

reg [5:0] mem_MUX [0:63];

always @* begin
  case (rot_mode)
    2'b00: begin
      for (i = 0; i < 64; i = i + 1)
        mem_MUX[i] = mem[i ^ 6'd0]; 
    end
    2'b01: begin
      for (i = 0; i < 64; i = i + 1)
        mem_MUX[i] = mem[i ^ 6'd1]; 
    end
    2'b10: begin
      for (i = 0; i < 64; i = i + 1)
        mem_MUX[i] = mem[i ^ 6'd2];
    end
    2'b11: begin
      for (i = 0; i < 64; i = i + 1)
        mem_MUX[i] = mem[i ^ 6'd3]; 
    end
    default: begin
      for (i = 0; i < 64; i = i + 1)
        mem_MUX[i] = mem[i];
    end
  endcase
end




always @(posedge clk) begin
	if (load) begin
		mem[63] <= rotorB_sram_din;
		for (i = 0; i < 63; i = i + 1)
			mem[i] <= mem[i+1];
	end
	else if (rotorB_in_valid) begin
		mem[0]  <= mem_MUX[56];
		mem[1]  <= mem_MUX[61];
		mem[2]  <= mem_MUX[25];
		mem[3]  <= mem_MUX[17];
		mem[4]  <= mem_MUX[42];
		mem[5]  <= mem_MUX[48];
		mem[6]  <= mem_MUX[23];
		mem[7]  <= mem_MUX[43];
		mem[8]  <= mem_MUX[10];
		mem[9]  <= mem_MUX[28];
		mem[10] <= mem_MUX[58];
		mem[11] <= mem_MUX[24];
		mem[12] <= mem_MUX[21];
		mem[13] <= mem_MUX[29];
		mem[14] <= mem_MUX[18];
		mem[15] <= mem_MUX[38];
		mem[16] <= mem_MUX[26];
		mem[17] <= mem_MUX[13];
		mem[18] <= mem_MUX[57];
		mem[19] <= mem_MUX[6];
		mem[20] <= mem_MUX[22];
		mem[21] <= mem_MUX[47];
		mem[22] <= mem_MUX[8];
		mem[23] <= mem_MUX[40];
		mem[24] <= mem_MUX[54];
		mem[25] <= mem_MUX[2];
		mem[26] <= mem_MUX[32];
		mem[27] <= mem_MUX[63];
		mem[28] <= mem_MUX[14];
		mem[29] <= mem_MUX[34];
		mem[30] <= mem_MUX[60];
		mem[31] <= mem_MUX[55];
		mem[32] <= mem_MUX[49];
		mem[33] <= mem_MUX[16];
		mem[34] <= mem_MUX[9];
		mem[35] <= mem_MUX[44];
		mem[36] <= mem_MUX[5];
		mem[37] <= mem_MUX[3];
		mem[38] <= mem_MUX[53];
		mem[39] <= mem_MUX[46];
		mem[40] <= mem_MUX[51];
		mem[41] <= mem_MUX[39];
		mem[42] <= mem_MUX[30];
		mem[43] <= mem_MUX[11];
		mem[44] <= mem_MUX[15];
		mem[45] <= mem_MUX[4];
		mem[46] <= mem_MUX[36];
		mem[47] <= mem_MUX[59];
		mem[48] <= mem_MUX[50];
		mem[49] <= mem_MUX[19];
		mem[50] <= mem_MUX[35];
		mem[51] <= mem_MUX[52];
		mem[52] <= mem_MUX[62];
		mem[53] <= mem_MUX[1];
		mem[54] <= mem_MUX[37];
		mem[55] <= mem_MUX[7];
		mem[56] <= mem_MUX[12];
		mem[57] <= mem_MUX[45];
		mem[58] <= mem_MUX[31];
		mem[59] <= mem_MUX[27];
		mem[60] <= mem_MUX[41];
		mem[61] <= mem_MUX[20];
		mem[62] <= mem_MUX[0];
		mem[63] <= mem_MUX[33];
	end
end

assign rotorB_for_dout = mem[rotorB_for_addr];




// for inverse searching
reg [63:0] hit;
integer k;

always @* begin
  for (k = 0; k < 64; k = k + 1) hit[k] = (rotorB_inv_din == mem[k]);
end

/*
always @* begin
  rotorB_inv_dout = 6'd0; // default to avoid latch
  case (rotorB_inv_din) // synopsys parallel_case full_case
    mem[0]  : rotorB_inv_dout = 6'd0;
    mem[1]  : rotorB_inv_dout = 6'd1;
    mem[2]  : rotorB_inv_dout = 6'd2;
    mem[3]  : rotorB_inv_dout = 6'd3;
    mem[4]  : rotorB_inv_dout = 6'd4;
    mem[5]  : rotorB_inv_dout = 6'd5;
    mem[6]  : rotorB_inv_dout = 6'd6;
    mem[7]  : rotorB_inv_dout = 6'd7;
    mem[8]  : rotorB_inv_dout = 6'd8;
    mem[9]  : rotorB_inv_dout = 6'd9;
    mem[10] : rotorB_inv_dout = 6'd10;
    mem[11] : rotorB_inv_dout = 6'd11;
    mem[12] : rotorB_inv_dout = 6'd12;
    mem[13] : rotorB_inv_dout = 6'd13;
    mem[14] : rotorB_inv_dout = 6'd14;
    mem[15] : rotorB_inv_dout = 6'd15;
    mem[16] : rotorB_inv_dout = 6'd16;
    mem[17] : rotorB_inv_dout = 6'd17;
    mem[18] : rotorB_inv_dout = 6'd18;
    mem[19] : rotorB_inv_dout = 6'd19;
    mem[20] : rotorB_inv_dout = 6'd20;
    mem[21] : rotorB_inv_dout = 6'd21;
    mem[22] : rotorB_inv_dout = 6'd22;
    mem[23] : rotorB_inv_dout = 6'd23;
    mem[24] : rotorB_inv_dout = 6'd24;
    mem[25] : rotorB_inv_dout = 6'd25;
    mem[26] : rotorB_inv_dout = 6'd26;
    mem[27] : rotorB_inv_dout = 6'd27;
    mem[28] : rotorB_inv_dout = 6'd28;
    mem[29] : rotorB_inv_dout = 6'd29;
    mem[30] : rotorB_inv_dout = 6'd30;
    mem[31] : rotorB_inv_dout = 6'd31;
    mem[32] : rotorB_inv_dout = 6'd32;
    mem[33] : rotorB_inv_dout = 6'd33;
    mem[34] : rotorB_inv_dout = 6'd34;
    mem[35] : rotorB_inv_dout = 6'd35;
    mem[36] : rotorB_inv_dout = 6'd36;
    mem[37] : rotorB_inv_dout = 6'd37;
    mem[38] : rotorB_inv_dout = 6'd38;
    mem[39] : rotorB_inv_dout = 6'd39;
    mem[40] : rotorB_inv_dout = 6'd40;
    mem[41] : rotorB_inv_dout = 6'd41;
    mem[42] : rotorB_inv_dout = 6'd42;
    mem[43] : rotorB_inv_dout = 6'd43;
    mem[44] : rotorB_inv_dout = 6'd44;
    mem[45] : rotorB_inv_dout = 6'd45;
    mem[46] : rotorB_inv_dout = 6'd46;
    mem[47] : rotorB_inv_dout = 6'd47;
    mem[48] : rotorB_inv_dout = 6'd48;
    mem[49] : rotorB_inv_dout = 6'd49;
    mem[50] : rotorB_inv_dout = 6'd50;
    mem[51] : rotorB_inv_dout = 6'd51;
    mem[52] : rotorB_inv_dout = 6'd52;
    mem[53] : rotorB_inv_dout = 6'd53;
    mem[54] : rotorB_inv_dout = 6'd54;
    mem[55] : rotorB_inv_dout = 6'd55;
    mem[56] : rotorB_inv_dout = 6'd56;
    mem[57] : rotorB_inv_dout = 6'd57;
    mem[58] : rotorB_inv_dout = 6'd58;
    mem[59] : rotorB_inv_dout = 6'd59;
    mem[60] : rotorB_inv_dout = 6'd60;
    mem[61] : rotorB_inv_dout = 6'd61;
    mem[62] : rotorB_inv_dout = 6'd62;
    mem[63] : rotorB_inv_dout = 6'd63;
    default : rotorB_inv_dout = 6'd0;
  endcase
end
*/


always @* begin
  rotorB_inv_dout = 6'd0;
  
  casez (hit) // synopsys parallel_case
    64'b???????????????????????????????????????????????????????????????1: rotorB_inv_dout = 6'd0;
    64'b??????????????????????????????????????????????????????????????1?: rotorB_inv_dout = 6'd1;
    64'b?????????????????????????????????????????????????????????????1??: rotorB_inv_dout = 6'd2;
    64'b????????????????????????????????????????????????????????????1???: rotorB_inv_dout = 6'd3;
    64'b???????????????????????????????????????????????????????????1????: rotorB_inv_dout = 6'd4;
    64'b??????????????????????????????????????????????????????????1?????: rotorB_inv_dout = 6'd5;
    64'b?????????????????????????????????????????????????????????1??????: rotorB_inv_dout = 6'd6;
    64'b????????????????????????????????????????????????????????1???????: rotorB_inv_dout = 6'd7;
    64'b???????????????????????????????????????????????????????1????????: rotorB_inv_dout = 6'd8;
    64'b??????????????????????????????????????????????????????1?????????: rotorB_inv_dout = 6'd9;
    64'b?????????????????????????????????????????????????????1??????????: rotorB_inv_dout = 6'd10;
    64'b????????????????????????????????????????????????????1???????????: rotorB_inv_dout = 6'd11;
    64'b???????????????????????????????????????????????????1????????????: rotorB_inv_dout = 6'd12;
    64'b??????????????????????????????????????????????????1?????????????: rotorB_inv_dout = 6'd13;
    64'b?????????????????????????????????????????????????1??????????????: rotorB_inv_dout = 6'd14;
    64'b????????????????????????????????????????????????1???????????????: rotorB_inv_dout = 6'd15;
    64'b???????????????????????????????????????????????1????????????????: rotorB_inv_dout = 6'd16;
    64'b??????????????????????????????????????????????1?????????????????: rotorB_inv_dout = 6'd17;
    64'b?????????????????????????????????????????????1??????????????????: rotorB_inv_dout = 6'd18;
    64'b????????????????????????????????????????????1???????????????????: rotorB_inv_dout = 6'd19;
    64'b???????????????????????????????????????????1????????????????????: rotorB_inv_dout = 6'd20;
    64'b??????????????????????????????????????????1?????????????????????: rotorB_inv_dout = 6'd21;
    64'b?????????????????????????????????????????1??????????????????????: rotorB_inv_dout = 6'd22;
    64'b????????????????????????????????????????1???????????????????????: rotorB_inv_dout = 6'd23;
    64'b???????????????????????????????????????1????????????????????????: rotorB_inv_dout = 6'd24;
    64'b??????????????????????????????????????1?????????????????????????: rotorB_inv_dout = 6'd25;
    64'b?????????????????????????????????????1??????????????????????????: rotorB_inv_dout = 6'd26;
    64'b????????????????????????????????????1???????????????????????????: rotorB_inv_dout = 6'd27;
    64'b???????????????????????????????????1????????????????????????????: rotorB_inv_dout = 6'd28;
    64'b??????????????????????????????????1?????????????????????????????: rotorB_inv_dout = 6'd29;
    64'b?????????????????????????????????1??????????????????????????????: rotorB_inv_dout = 6'd30;
    64'b????????????????????????????????1???????????????????????????????: rotorB_inv_dout = 6'd31;
    64'b???????????????????????????????1????????????????????????????????: rotorB_inv_dout = 6'd32;
    64'b??????????????????????????????1?????????????????????????????????: rotorB_inv_dout = 6'd33;
    64'b?????????????????????????????1??????????????????????????????????: rotorB_inv_dout = 6'd34;
    64'b????????????????????????????1???????????????????????????????????: rotorB_inv_dout = 6'd35;
    64'b???????????????????????????1????????????????????????????????????: rotorB_inv_dout = 6'd36;
    64'b??????????????????????????1?????????????????????????????????????: rotorB_inv_dout = 6'd37;
    64'b?????????????????????????1??????????????????????????????????????: rotorB_inv_dout = 6'd38;
    64'b????????????????????????1???????????????????????????????????????: rotorB_inv_dout = 6'd39;
    64'b???????????????????????1????????????????????????????????????????: rotorB_inv_dout = 6'd40;
    64'b??????????????????????1?????????????????????????????????????????: rotorB_inv_dout = 6'd41;
    64'b?????????????????????1??????????????????????????????????????????: rotorB_inv_dout = 6'd42;
    64'b????????????????????1???????????????????????????????????????????: rotorB_inv_dout = 6'd43;
    64'b???????????????????1????????????????????????????????????????????: rotorB_inv_dout = 6'd44;
    64'b??????????????????1?????????????????????????????????????????????: rotorB_inv_dout = 6'd45;
    64'b?????????????????1??????????????????????????????????????????????: rotorB_inv_dout = 6'd46;
    64'b????????????????1???????????????????????????????????????????????: rotorB_inv_dout = 6'd47;
    64'b???????????????1????????????????????????????????????????????????: rotorB_inv_dout = 6'd48;
    64'b??????????????1?????????????????????????????????????????????????: rotorB_inv_dout = 6'd49;
    64'b?????????????1??????????????????????????????????????????????????: rotorB_inv_dout = 6'd50;
    64'b????????????1???????????????????????????????????????????????????: rotorB_inv_dout = 6'd51;
    64'b???????????1????????????????????????????????????????????????????: rotorB_inv_dout = 6'd52;
    64'b??????????1?????????????????????????????????????????????????????: rotorB_inv_dout = 6'd53;
    64'b?????????1??????????????????????????????????????????????????????: rotorB_inv_dout = 6'd54;
    64'b????????1???????????????????????????????????????????????????????: rotorB_inv_dout = 6'd55;
    64'b???????1????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd56;
    64'b??????1?????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd57;
    64'b?????1??????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd58;
    64'b????1???????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd59;
    64'b???1????????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd60;
    64'b??1?????????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd61;
    64'b?1??????????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd62;
    64'b1???????????????????????????????????????????????????????????????: rotorB_inv_dout = 6'd63;
    default: ; 
  endcase
end


endmodule

module inverse_mapping (
  input [1:0] mode,
  input [5:0] din,
  output reg [5:0] dout
);

wire [5:0] xor_din;

assign xor_din = din ^ {4'd0, mode};

always @* begin
  case (xor_din)
    6'h00: dout = 6'h38; // 56
    6'h01: dout = 6'h3D; // 61
    6'h02: dout = 6'h19; // 25
    6'h03: dout = 6'h11; // 17
    6'h04: dout = 6'h2A; // 42
    6'h05: dout = 6'h30; // 48
    6'h06: dout = 6'h17; // 23
    6'h07: dout = 6'h2B; // 43
    6'h08: dout = 6'h0A; // 10
    6'h09: dout = 6'h1C; // 28
    6'h0A: dout = 6'h3A; // 58
    6'h0B: dout = 6'h18; // 24
    6'h0C: dout = 6'h15; // 21
    6'h0D: dout = 6'h1D; // 29
    6'h0E: dout = 6'h12; // 18
    6'h0F: dout = 6'h26; // 38
    6'h10: dout = 6'h1A; // 26
    6'h11: dout = 6'h0D; // 13
    6'h12: dout = 6'h39; // 57
    6'h13: dout = 6'h06; // 06
    6'h14: dout = 6'h16; // 22
    6'h15: dout = 6'h2F; // 47
    6'h16: dout = 6'h08; // 08
    6'h17: dout = 6'h28; // 40
    6'h18: dout = 6'h36; // 54
    6'h19: dout = 6'h02; // 02
    6'h1A: dout = 6'h20; // 32
    6'h1B: dout = 6'h3F; // 63
    6'h1C: dout = 6'h0E; // 14
    6'h1D: dout = 6'h22; // 34
    6'h1E: dout = 6'h3C; // 60
    6'h1F: dout = 6'h37; // 55
    6'h20: dout = 6'h31; // 49
    6'h21: dout = 6'h10; // 16
    6'h22: dout = 6'h09; // 09
    6'h23: dout = 6'h2C; // 44
    6'h24: dout = 6'h05; // 05
    6'h25: dout = 6'h03; // 03
    6'h26: dout = 6'h35; // 53
    6'h27: dout = 6'h2E; // 46
    6'h28: dout = 6'h33; // 51
    6'h29: dout = 6'h27; // 39
    6'h2A: dout = 6'h1E; // 30
    6'h2B: dout = 6'h0B; // 11
    6'h2C: dout = 6'h0F; // 15
    6'h2D: dout = 6'h04; // 04
    6'h2E: dout = 6'h24; // 36
    6'h2F: dout = 6'h3B; // 59
    6'h30: dout = 6'h32; // 50
    6'h31: dout = 6'h13; // 19
    6'h32: dout = 6'h23; // 35
    6'h33: dout = 6'h34; // 52
    6'h34: dout = 6'h3E; // 62
    6'h35: dout = 6'h01; // 01
    6'h36: dout = 6'h25; // 37
    6'h37: dout = 6'h07; // 07
    6'h38: dout = 6'h0C; // 12
    6'h39: dout = 6'h2D; // 45
    6'h3A: dout = 6'h1F; // 31
    6'h3B: dout = 6'h1B; // 27
    6'h3C: dout = 6'h29; // 41
    6'h3D: dout = 6'h14; // 20
    6'h3E: dout = 6'h00; // 00
    6'h3F: dout = 6'h21; // 33
    default: dout = 6'h00;
  endcase
end


endmodule